`define DATA_WIDTH 9

`define FIFO_PTR_WIDTH 4
`define FIFO_DEPTH 16
`define FIFO_FULL_BIT 4
`define PTR_WIDTH 3

`define PACKET_LEN_MSB 7
`define PACKET_LEN_LSB 2
